-- Add your stimulus here ...
process
begin
x <= "0000000000000111";
y <= "0000000000010000";
Cin <= '0';
wait for 10 ns;
x <= "0000000000001111";
y <= "0000000000010000";
Cin <= '0';
wait for 10 ns;
x <= "0000000001000111";
y <= "0000000000011000";
Cin <= '0';
wait for 10 ns;
x <= "0000001110000111";
y <= "0000000110010000";
Cin <= '0';
wait for 10 ns;
x <= "0000000000110111";
y <= "0000001100010000";
Cin <= '0';
wait for 10 ns;
x <= "0000000100000111";
y <= "0000000000110000";
Cin <= '0';
wait for 10 ns;
x <= "0000000000100111";
y <= "0001000000010000";
Cin <= '0';
wait for 10 ns;
end process;
